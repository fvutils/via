
typedef class via_object_type_if;

class via_object_if;

    virtual function via_object_type_if get_object_type();
    endfunction

endclass

