
typedef class via_visitor;

interface class via_accept_if;

    pure virtual function void accept(via_visitor v);

endclass