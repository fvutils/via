
typedef class via_visitor;

class via_accept_if;

    virtual function void accept(via_visitor v);
    endfunction

endclass