
// Defines the interface between an environment and its roots
class via_root_if;

endclass