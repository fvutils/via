
class via_component_if;

    virtual function string get_name();
    endfunction

    virtual function string get_full_name();
    endfunction
endclass
