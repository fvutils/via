
typedef class via_field;

class via_object_type_if;
    via_field fields[$];

    virtual function string get_name();
    endfunction

    virtual function void get_fields(via_field fields[$]);
    endfunction

endclass
