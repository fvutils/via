


class via_uvm_classtype_factory;


endclass
