

class via_analysis_port_subscriber;

    virtual function void write(via_object t);
    endfunction

endclass
