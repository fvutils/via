
typedef interface class via_component_if;

interface class via_sequencer_if extends via_component_if;

endclass

