
`ifndef INCLUDED_VIA_MACROS_SVH
`define INCLUDED_VIA_MACROS_SVH

`endif /* INCLUDED_VIA_MACROS_SVH */

