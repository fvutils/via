
package via;

    `include "via_component_if.svh"
    `include "via_root.svh"
    `include "via_root_listener_if.svh"

endpackage

