
class via_analysis_port_if;

    virtual function void add_listener(via_analysis_port_listener l);
    endfunction

endclass
