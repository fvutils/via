
interface class via_factory_if;

    pure virtual function void get_type_names(ref string names[$]);

endclass