
class via_uvm_object extends via_object_if;
    uvm_object      obj;


endclass
