
package test_utils;
    import via::*;

    `include "type_finder.svh"

endpackage

