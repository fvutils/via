
typedef class via_field;

class via_class_type;
    string name;
    via_field fields[$];

    function new(string name);
        this.name = name;
    endfunction

endclass
